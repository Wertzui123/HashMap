module hashmap

fn modulo(a int, b int) int {
	return ((a % b) + b) % b
}
